module Instruction_Mem(
	input		[31:0]	PC_F,
	input			clk,
	input			rst,
	output	reg	[31:0]	instruction
);

reg	[31:0]	instrmem [16:0];

always @(posedge clk or posedge rst) begin
	if(rst) begin
		instruction	<= 0;
		instrmem[0]	<= 32'b100100_00000_00000_01001_0001_0001_001;
		instrmem[1]	<= 32'b100100_00000_00000_01010_0001_0001_001;
		instrmem[2]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[3]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[4]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[5]	<= 32'b100001_00000_01001_00000_0000_0000_000;
		instrmem[6]	<= 32'b110000_01001_01010_01011_00000_000001;
		instrmem[7]	<= 32'b100000_00000_00000_01101_00000_000000;
		instrmem[8]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[9]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[10]	<= 32'b000000_00000_00000_00000_0000_0000_000;
		instrmem[11]	<= 32'b010101_01101_01001_01100_00000_100001;
		instrmem[12] 	<= 0;
		instrmem[13]	<= 0;
		instrmem[14]	<= 0;
		instrmem[15]	<= 0;
	end
	
	else begin
		instruction <= instrmem[PC_F >> 2];
	end
end

/* initial begin
	$readmemb("instructions.txt", instrmem);
end */

/* initial begin
	instrmem[0]	= 32'b100100_00000_00000_01001_0001_0001_001;
	instrmem[1]	= 32'b100100_00000_00000_01010_0001_0001_001;
	instrmem[2]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[3]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[4]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[5]	= 32'b100001_00000_01001_00000_0000_0000_000;
	instrmem[6]	= 32'b110000_01001_01010_01011_00000_000001;
	instrmem[7]	= 32'b100000_00000_00000_01101_00000_000000;
	instrmem[8]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[9]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[10]	= 32'b000000_00000_00000_00000_0000_0000_000;
	instrmem[11]	= 32'b010101_01101_01001_01100_00000_100001;
end */

endmodule

